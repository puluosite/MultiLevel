** 40 cascaded, 2 paralleled cells


**First Colony Starts
**it does not exit, short!
R111_1 1 11_1 1e-30

**it does not exit, short!
R11_111_2 11_1 11_2 1e-30

I11_211_3 11_3 11_2_0 DC 3.000000e+00
D11_211_3 11_2_0 11_3 diode11_211_3
Rs11_211_3 11_2 11_2_0 4.740000e-02
Rsh11_211_3 11_2_0 11_3 5.000000e+03
.MODEL diode11_211_3 D IS=1.000000e-06 N=9.000000e+00

**it does not exit, short!
R11_311_4 11_3 11_4 1e-30

I11_411 11 11_4_0 DC 2.000000e+00
D11_411 11_4_0 11 diode11_411
Rs11_411 11_4 11_4_0 5.530000e-02
Rsh11_411 11_4_0 11 5.000000e+03
.MODEL diode11_411 D IS=1.000000e-06 N=1.050000e+01

.MODEL diode_bp111 D IS=1.000000e-05 N=1.000000e+00
D_Bypass111 11 1 diode_bp111

**Second Colony Starts
**it does not exit, short!
R1121_1 11 21_1 1e-30

I21_121_2 21_2 21_1_0 DC 3.500000e+00
D21_121_2 21_1_0 21_2 diode21_121_2
Rs21_121_2 21_1 21_1_0 3.950000e-02
Rsh21_121_2 21_1_0 21_2 5.000000e+03
.MODEL diode21_121_2 D IS=1.000000e-06 N=7.500000e+00

**it does not exit, short!
R21_221_3 21_2 21_3 1e-30

**it does not exit, short!
R21_321_4 21_3 21_4 1e-30

I21_421 21 21_4_0 DC 2.000000e+00
D21_421 21_4_0 21 diode21_421
Rs21_421 21_4 21_4_0 6.320000e-02
Rsh21_421 21_4_0 21 5.000000e+03
.MODEL diode21_421 D IS=1.000000e-06 N=1.200000e+01

.MODEL diode_bp2111 D IS=1.000000e-05 N=1.000000e+00
D_Bypass2111 21 11 diode_bp2111

**Third Colony Starts
I2131_1 31_1 21_0 DC 4.000000e+00
D2131_1 21_0 31_1 diode2131_1
Rs2131_1 21 21_0 1.027000e-01
Rsh2131_1 21_0 31_1 5.000000e+03
.MODEL diode2131_1 D IS=1.000000e-06 N=1.950000e+01

**it does not exit, short!
R31_131_2 31_1 31_2 1e-30

**it does not exit, short!
R31_231_3 31_2 31_3 1e-30

**it does not exit, short!
R31_331_4 31_3 31_4 1e-30

I31_40 0 31_4_0 DC 2.000000e+00
D31_40 31_4_0 0 diode31_40
Rs31_40 31_4 31_4_0 7.900000e-03
Rsh31_40 31_4_0 0 5.000000e+03
.MODEL diode31_40 D IS=1.000000e-06 N=1.500000e+00

.MODEL diode_bp021 D IS=1.000000e-05 N=1.000000e+00
D_Bypass021 0 21 diode_bp021

**First Colony Starts
**it does not exit, short!
R112_1 1 12_1 1e-30

**it does not exit, short!
R12_112_2 12_1 12_2 1e-30

I12_212_3 12_3 12_2_0 DC 3.000000e+00
D12_212_3 12_2_0 12_3 diode12_212_3
Rs12_212_3 12_2 12_2_0 4.740000e-02
Rsh12_212_3 12_2_0 12_3 5.000000e+03
.MODEL diode12_212_3 D IS=1.000000e-06 N=9.000000e+00

**it does not exit, short!
R12_312_4 12_3 12_4 1e-30

I12_412 12 12_4_0 DC 2.000000e+00
D12_412 12_4_0 12 diode12_412
Rs12_412 12_4 12_4_0 5.530000e-02
Rsh12_412 12_4_0 12 5.000000e+03
.MODEL diode12_412 D IS=1.000000e-06 N=1.050000e+01

.MODEL diode_bp121 D IS=1.000000e-05 N=1.000000e+00
D_Bypass121 12 1 diode_bp121

**Second Colony Starts
**it does not exit, short!
R1222_1 12 22_1 1e-30

I22_122_2 22_2 22_1_0 DC 3.500000e+00
D22_122_2 22_1_0 22_2 diode22_122_2
Rs22_122_2 22_1 22_1_0 4.740000e-02
Rsh22_122_2 22_1_0 22_2 5.000000e+03
.MODEL diode22_122_2 D IS=1.000000e-06 N=9.000000e+00

**it does not exit, short!
R22_222_3 22_2 22_3 1e-30

I22_322_4 22_4 22_3_0 DC 2.500000e+00
D22_322_4 22_3_0 22_4 diode22_322_4
Rs22_322_4 22_3 22_3_0 5.530000e-02
Rsh22_322_4 22_3_0 22_4 5.000000e+03
.MODEL diode22_322_4 D IS=1.000000e-06 N=1.050000e+01

**it does not exit, short!
R22_422 22_4 22 1e-30

.MODEL diode_bp2212 D IS=1.000000e-05 N=1.000000e+00
D_Bypass2212 22 12 diode_bp2212

**Third Colony Starts
I2232_1 32_1 22_0 DC 4.000000e+00
D2232_1 22_0 32_1 diode2232_1
Rs2232_1 22 22_0 9.480000e-02
Rsh2232_1 22_0 32_1 5.000000e+03
.MODEL diode2232_1 D IS=1.000000e-06 N=1.800000e+01

**it does not exit, short!
R32_132_2 32_1 32_2 1e-30

**it does not exit, short!
R32_232_3 32_2 32_3 1e-30

**it does not exit, short!
R32_332_4 32_3 32_4 1e-30

I32_40 0 32_4_0 DC 2.000000e+00
D32_40 32_4_0 0 diode32_40
Rs32_40 32_4 32_4_0 1.580000e-02
Rsh32_40 32_4_0 0 5.000000e+03
.MODEL diode32_40 D IS=1.000000e-06 N=3.000000e+00

.MODEL diode_bp022 D IS=1.000000e-05 N=1.000000e+00
D_Bypass022 0 22 diode_bp022



 Vds 1 0
.DC Vds 0 60.000000 0.005
.PRINT V(1) I(Vds)
.end
