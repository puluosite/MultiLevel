** 30 cascaded, 4 paralleled cells


** subcircuit:4.000000e+00A,unshaded
.SUBCKT CELL1 P M 
 I1 M Y DC 4.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:3.500000e+00A,unshaded
.SUBCKT CELL2 P M 
 I1 M Y DC 3.500000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:3.000000e+00A,unshaded
.SUBCKT CELL3 P M 
 I1 M Y DC 3.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:2.500000e+00A,unshaded
.SUBCKT CELL4 P M 
 I1 M Y DC 2.500000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:2.000000e+00A,unshaded
.SUBCKT CELL5 P M 
 I1 M Y DC 2.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


 XU11 1 11 CELL5
 XU21 11 21 CELL5
 XU31 21 31 CELL5
 XU41 31 41 CELL5
 XU51 41 51 CELL5
 XU61 51 61 CELL4
 XU71 61 71 CELL4
 XU81 71 81 CELL4
 XU91 81 91 CELL4
 XU101 91 101 CELL4
 XU111 101 111 CELL4
 XU121 111 121 CELL4
 XU131 121 131 CELL4
 XU141 131 141 CELL3
 XU151 141 151 CELL2
 XU161 151 161 CELL2
 XU171 161 171 CELL2
 XU181 171 181 CELL2
 XU191 181 191 CELL1
 XU201 191 201 CELL1
 XU211 201 211 CELL1
 XU221 211 221 CELL1
 XU231 221 231 CELL1
 XU241 231 241 CELL1
 XU251 241 251 CELL1
 XU261 251 261 CELL1
 XU271 261 271 CELL1
 XU281 271 281 CELL2
 XU291 281 291 CELL2
 XU301 291 0 CELL3

 D_Bypass11 0 151  diode_b1

 D_Bypass21 151 1  diode_b1
.MODEL diode_b1 D IS=1.000000e-05 N=1.000000e+00
 XU12 1 12 CELL5
 XU22 12 22 CELL5
 XU32 22 32 CELL5
 XU42 32 42 CELL5
 XU52 42 52 CELL5
 XU62 52 62 CELL5
 XU72 62 72 CELL4
 XU82 72 82 CELL4
 XU92 82 92 CELL4
 XU102 92 102 CELL4
 XU112 102 112 CELL4
 XU122 112 122 CELL3
 XU132 122 132 CELL3
 XU142 132 142 CELL2
 XU152 142 152 CELL2
 XU162 152 162 CELL2
 XU172 162 172 CELL2
 XU182 172 182 CELL1
 XU192 182 192 CELL1
 XU202 192 202 CELL1
 XU212 202 212 CELL1
 XU222 212 222 CELL2
 XU232 222 232 CELL1
 XU242 232 242 CELL1
 XU252 242 252 CELL1
 XU262 252 262 CELL1
 XU272 262 272 CELL1
 XU282 272 282 CELL1
 XU292 282 292 CELL2
 XU302 292 0 CELL3

 D_Bypass12 0 152  diode_b2

 D_Bypass22 152 1  diode_b2
.MODEL diode_b2 D IS=1.000000e-05 N=1.000000e+00
 XU13 1 13 CELL5
 XU23 13 23 CELL5
 XU33 23 33 CELL5
 XU43 33 43 CELL5
 XU53 43 53 CELL5
 XU63 53 63 CELL5
 XU73 63 73 CELL4
 XU83 73 83 CELL4
 XU93 83 93 CELL4
 XU103 93 103 CELL4
 XU113 103 113 CELL4
 XU123 113 123 CELL3
 XU133 123 133 CELL3
 XU143 133 143 CELL3
 XU153 143 153 CELL2
 XU163 153 163 CELL2
 XU173 163 173 CELL2
 XU183 173 183 CELL2
 XU193 183 193 CELL1
 XU203 193 203 CELL1
 XU213 203 213 CELL1
 XU223 213 223 CELL1
 XU233 223 233 CELL1
 XU243 233 243 CELL1
 XU253 243 253 CELL1
 XU263 253 263 CELL5
 XU273 263 273 CELL1
 XU283 273 283 CELL2
 XU293 283 293 CELL2
 XU303 293 0 CELL3

 D_Bypass13 0 153  diode_b3

 D_Bypass23 153 1  diode_b3
.MODEL diode_b3 D IS=1.000000e-05 N=1.000000e+00
 XU14 1 14 CELL5
 XU24 14 24 CELL5
 XU34 24 34 CELL5
 XU44 34 44 CELL5
 XU54 44 54 CELL5
 XU64 54 64 CELL5
 XU74 64 74 CELL4
 XU84 74 84 CELL4
 XU94 84 94 CELL4
 XU104 94 104 CELL4
 XU114 104 114 CELL4
 XU124 114 124 CELL4
 XU134 124 134 CELL3
 XU144 134 144 CELL3
 XU154 144 154 CELL2
 XU164 154 164 CELL2
 XU174 164 174 CELL2
 XU184 174 184 CELL2
 XU194 184 194 CELL1
 XU204 194 204 CELL1
 XU214 204 214 CELL1
 XU224 214 224 CELL1
 XU234 224 234 CELL1
 XU244 234 244 CELL1
 XU254 244 254 CELL1
 XU264 254 264 CELL1
 XU274 264 274 CELL1
 XU284 274 284 CELL2
 XU294 284 294 CELL2
 XU304 294 0 CELL3

 D_Bypass14 0 154  diode_b4

 D_Bypass24 154 1  diode_b4
.MODEL diode_b4 D IS=1.000000e-05 N=1.000000e+00


 Vds 1 0
.DC Vds 0 30.000000 0.005
.PRINT V(1) I(Vds)
.end
