** 60 cascaded, 2 paralleled cells


** subcircuit:4.000000e+00A,unshaded
.SUBCKT CELL1 P M 
 I1 M Y DC 4.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:3.500000e+00A,unshaded
.SUBCKT CELL2 P M 
 I1 M Y DC 3.500000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:3.000000e+00A,unshaded
.SUBCKT CELL3 P M 
 I1 M Y DC 3.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:2.500000e+00A,unshaded
.SUBCKT CELL4 P M 
 I1 M Y DC 2.500000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:2.000000e+00A,unshaded
.SUBCKT CELL5 P M 
 I1 M Y DC 2.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


 XU11 1 11 CELL5
 XU21 11 21 CELL5
 XU31 21 31 CELL5
 XU41 31 41 CELL5
 XU51 41 51 CELL5
 XU61 51 61 CELL4
 XU71 61 71 CELL4
 XU81 71 81 CELL4
 XU91 81 91 CELL5
 XU101 91 101 CELL3
 XU111 101 111 CELL4
 XU121 111 121 CELL3
 XU131 121 131 CELL2
 XU141 131 141 CELL2
 XU151 141 151 CELL2
 XU161 151 161 CELL2
 XU171 161 171 CELL2
 XU181 171 181 CELL1
 XU191 181 191 CELL1
 XU201 191 201 CELL1
 XU211 201 211 CELL1
 XU221 211 221 CELL1
 XU231 221 231 CELL1
 XU241 231 241 CELL1
 XU251 241 251 CELL1
 XU261 251 261 CELL1
 XU271 261 271 CELL1
 XU281 271 281 CELL1
 XU291 281 291 CELL1
 XU301 291 301 CELL1
 XU311 301 311 CELL1
 XU321 311 321 CELL1
 XU331 321 331 CELL1
 XU341 331 341 CELL1
 XU351 341 351 CELL1
 XU361 351 361 CELL1
 XU371 361 371 CELL1
 XU381 371 381 CELL1
 XU391 381 391 CELL1
 XU401 391 401 CELL1
 XU411 401 411 CELL1
 XU421 411 421 CELL1
 XU431 421 431 CELL1
 XU441 431 441 CELL1
 XU451 441 451 CELL1
 XU461 451 461 CELL1
 XU471 461 471 CELL1
 XU481 471 481 CELL1
 XU491 481 491 CELL1
 XU501 491 501 CELL1
 XU511 501 511 CELL1
 XU521 511 521 CELL1
 XU531 521 531 CELL1
 XU541 531 541 CELL1
 XU551 541 551 CELL1
 XU561 551 561 CELL1
 XU571 561 571 CELL1
 XU581 571 581 CELL1
 XU591 581 591 CELL1
 XU601 591 0 CELL1

 D_Bypass11 0 401  diode_b1

 D_Bypass21 401 201  diode_b1

 D_Bypass31 201 1  diode_b1
.MODEL diode_b1 D IS=1.000000e-05 N=1.000000e+00
 XU12 1 12 CELL5
 XU22 12 22 CELL5
 XU32 22 32 CELL5
 XU42 32 42 CELL5
 XU52 42 52 CELL5
 XU62 52 62 CELL5
 XU72 62 72 CELL4
 XU82 72 82 CELL4
 XU92 82 92 CELL3
 XU102 92 102 CELL3
 XU112 102 112 CELL3
 XU122 112 122 CELL2
 XU132 122 132 CELL2
 XU142 132 142 CELL2
 XU152 142 152 CELL2
 XU162 152 162 CELL2
 XU172 162 172 CELL2
 XU182 172 182 CELL1
 XU192 182 192 CELL1
 XU202 192 202 CELL1
 XU212 202 212 CELL1
 XU222 212 222 CELL1
 XU232 222 232 CELL1
 XU242 232 242 CELL1
 XU252 242 252 CELL1
 XU262 252 262 CELL1
 XU272 262 272 CELL1
 XU282 272 282 CELL1
 XU292 282 292 CELL1
 XU302 292 302 CELL1
 XU312 302 312 CELL1
 XU322 312 322 CELL1
 XU332 322 332 CELL1
 XU342 332 342 CELL1
 XU352 342 352 CELL1
 XU362 352 362 CELL1
 XU372 362 372 CELL1
 XU382 372 382 CELL1
 XU392 382 392 CELL1
 XU402 392 402 CELL1
 XU412 402 412 CELL1
 XU422 412 422 CELL1
 XU432 422 432 CELL1
 XU442 432 442 CELL1
 XU452 442 452 CELL1
 XU462 452 462 CELL1
 XU472 462 472 CELL1
 XU482 472 482 CELL3
 XU492 482 492 CELL1
 XU502 492 502 CELL1
 XU512 502 512 CELL1
 XU522 512 522 CELL1
 XU532 522 532 CELL1
 XU542 532 542 CELL1
 XU552 542 552 CELL1
 XU562 552 562 CELL1
 XU572 562 572 CELL1
 XU582 572 582 CELL1
 XU592 582 592 CELL1
 XU602 592 0 CELL2

 D_Bypass12 0 402  diode_b2

 D_Bypass22 402 202  diode_b2

 D_Bypass32 202 1  diode_b2
.MODEL diode_b2 D IS=1.000000e-05 N=1.000000e+00


 Vds 1 0
.DC Vds 0 60.000000 0.005
.PRINT V(1) I(Vds)
.end
