** 40 cascaded, 2 paralleled cells


** subcircuit:4.000000e+00A,unshaded
.SUBCKT CELL1 P M 
 I1 M Y DC 4.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:3.500000e+00A,unshaded
.SUBCKT CELL2 P M 
 I1 M Y DC 3.500000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:3.000000e+00A,unshaded
.SUBCKT CELL3 P M 
 I1 M Y DC 3.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:2.500000e+00A,unshaded
.SUBCKT CELL4 P M 
 I1 M Y DC 2.500000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


** subcircuit:2.000000e+00A,unshaded
.SUBCKT CELL5 P M 
 I1 M Y DC 2.000000e+00
 D1 Y M diode1
 Rsh Y M 5.000000e+03
 Rs Y P 7.900000e-03
.MODEL diode1 D IS=1.000000e-06 N=1.500000e+00
.ENDS


 XU11 1 11 CELL5
 XU21 11 21 CELL5
 XU31 21 31 CELL5
 XU41 31 41 CELL5
 XU51 41 51 CELL5
 XU61 51 61 CELL5
 XU71 61 71 CELL4
 XU81 71 81 CELL3
 XU91 81 91 CELL3
 XU101 91 101 CELL3
 XU111 101 111 CELL3
 XU121 111 121 CELL3
 XU131 121 131 CELL3
 XU141 131 141 CELL3
 XU151 141 151 CELL3
 XU161 151 161 CELL4
 XU171 161 171 CELL4
 XU181 171 181 CELL4
 XU191 181 191 CELL4
 XU201 191 201 CELL4
 XU211 201 211 CELL4
 XU221 211 221 CELL4
 XU231 221 231 CELL5
 XU241 231 241 CELL2
 XU251 241 251 CELL2
 XU261 251 261 CELL2
 XU271 261 271 CELL2
 XU281 271 281 CELL2
 XU291 281 291 CELL2
 XU301 291 301 CELL2
 XU311 301 311 CELL5
 XU321 311 321 CELL1
 XU331 321 331 CELL1
 XU341 331 341 CELL1
 XU351 341 351 CELL1
 XU361 351 361 CELL1
 XU371 361 371 CELL1
 XU381 371 381 CELL1
 XU391 381 391 CELL1
 XU401 391 0 CELL1

 D_Bypass11 0 261  diode_b1

 D_Bypass21 261 131  diode_b1

 D_Bypass31 131 1  diode_b1
.MODEL diode_b1 D IS=1.000000e-05 N=1.000000e+00
 XU12 1 12 CELL5
 XU22 12 22 CELL5
 XU32 22 32 CELL5
 XU42 32 42 CELL5
 XU52 42 52 CELL5
 XU62 52 62 CELL5
 XU72 62 72 CELL4
 XU82 72 82 CELL3
 XU92 82 92 CELL3
 XU102 92 102 CELL3
 XU112 102 112 CELL3
 XU122 112 122 CELL3
 XU132 122 132 CELL3
 XU142 132 142 CELL3
 XU152 142 152 CELL4
 XU162 152 162 CELL3
 XU172 162 172 CELL4
 XU182 172 182 CELL4
 XU192 182 192 CELL4
 XU202 192 202 CELL4
 XU212 202 212 CELL4
 XU222 212 222 CELL4
 XU232 222 232 CELL2
 XU242 232 242 CELL2
 XU252 242 252 CELL2
 XU262 252 262 CELL2
 XU272 262 272 CELL2
 XU282 272 282 CELL2
 XU292 282 292 CELL2
 XU302 292 302 CELL2
 XU312 302 312 CELL2
 XU322 312 322 CELL5
 XU332 322 332 CELL1
 XU342 332 342 CELL1
 XU352 342 352 CELL1
 XU362 352 362 CELL1
 XU372 362 372 CELL1
 XU382 372 382 CELL1
 XU392 382 392 CELL1
 XU402 392 0 CELL5

 D_Bypass12 0 262  diode_b2

 D_Bypass22 262 132  diode_b2

 D_Bypass32 132 1  diode_b2
.MODEL diode_b2 D IS=1.000000e-05 N=1.000000e+00


 Vds 1 0
.DC Vds 0 60.000000 0.005
.PRINT V(1) I(Vds)
.end
